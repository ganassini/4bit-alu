LIBRARY	IEEE;
USE IEEE.std_logic_1164.all;

ENTITY seg7 IS
  PORT(
    entrada: IN std_logic_vector(3 downto 0);
    zero: OUT std_logic_vector(0 downto 0);
    s: OUT std_logic_vector(41 downto 0)
  );
END seg7;

ARCHITECTURE arq_seg7 OF seg7 IS
BEGIN 
  with entrada select
    s <= "100000010000001000000100000010000001000000" when "0000",
         "100000011110011000000100000010000001111001" when "0001",
     	 "100000001001001000000100000011110011000000" when "0010",
         "100000001100001000000100000011110011111001" when "0011",
         "100000000110011000000111100110000001000000" when "0100",
         "100000000100101000000111100110000001111001" when "0101",
         "100000000000101000000111100111110011000000" when "0110",
         "100000011110001000000111100111110011111001" when "0111",
         "100000000000001111001100000010000001000000" when "1000",
         "100000000100001111001100000010000001111001" when "1001",
         "111100110000001111001100000011110011000000" when "1010",
         "111100111110011111001100000011110011111001" when "1011",
         "111100101001001111001111100110000001000000" when "1100",
         "111100101100001111001111100110000001111001" when "1101",
         "111100100110011111001111100111110011000000" when "1110",
         "111100100100101111001111100111110011111001" when "1111",
         "011111101111110111111011111101111110111111" when others;
 
  with entrada select
    zero <= "1" when "0000",
      	    "0" when others;  
END arq_seg7;
